class alu_generator;

rand alu_transaction trans;
